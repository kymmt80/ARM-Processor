module EXE_stage (
    input clk,rst,
    input[31:0] PC_in,
    output [31:0] PC
);
endmodule


module EXE_Stage_Reg (
    input clk,rst,
    input[31:0] PC_in,
    output [31:0] PC
);
endmodule