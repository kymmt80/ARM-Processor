module MEM_stage (
    input clk,rst,
    input[31:0] PC_in,
    output [31:0] PC
);
endmodule


module MEM_Stage_Reg (
    input clk,rst,
    input[31:0] PC_in,
    output [31:0] PC
);
endmodule