module data_mem(input memWrite,memRead,input [31:0]writeData,Address,output reg [31:0]readData);
reg[31:0] mem[0:65535];

initial begin
    mem[1000]=32'b11111111111111111111111110011100;
    mem[1004]=32'b00000000000000000000000000000000;
    mem[1008]=32'b00000000000000000000000000000101;
    mem[1012]=32'b00000000000000000000000000000101;
    mem[1016]=32'b00000000000000000000000000000101;
    mem[1020]=32'b00000000000000000000000000000101;
    mem[1024]=32'b11111111111111111111111101101010;
    mem[1028]=32'b00000000000000000000000000000000;
    mem[1032]=32'b00000000000000000000000000000001;
    mem[1036]=32'b00000000000000000000000000000001;
end

always@(memRead,Address)begin
    if (memRead ==1)
        readData <= mem[((Address>>2)<<2)-32'd1024];
end

always@(posedge clk)begin
    if(memWrite==1)
        mem[((Address>>2)<<2)-32'd1024]<=writeData;
end
endmodule