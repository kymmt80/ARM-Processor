module hazard_Detection_unit(
    input [3:0]src1,
    input [3:0]src2,
    input [3:0]Exe_Dest,
    input Exe_WB_EN,
    input [3:0]Mem_Dest,
    input Mem_WB_EN,
    output hazard_Detected);

endmodule