module ID_stage (
    input clk,rst,
    input[31:0] PC_in,
    output [31:0] PC
);
endmodule


module ID_Stage_Reg (
    input clk,rst,
    input[31:0] PC_in,
    output [31:0] PC
);
endmodule