module Condition_Check(
    input Cond,
    input[3:0] SR,
    output check_output);
endmodule