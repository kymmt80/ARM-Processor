module inst_mem(input [31:0]Address,output reg [31:0]inst);
reg [31:0] mem[0:127];

initial begin
    
mem[1-1]=32'b1110_00_1_1101_0_0000_0000_000000010100; //MOV		R0 ,#20 		//R0 = 20
mem[2-1]=32'b1110_00_1_1101_0_0000_0001_101000000001; //MOV		R1 ,#4096		//R1 = 4096
mem[3-1]=32'b1110_00_1_1101_0_0000_0010_000100000011; //MOV		R2 ,#0xC0000000	//R2 = -1073741824
mem[4-1]=32'b1110_00_0_0100_1_0010_0011_000000000010; //ADDS		R3 ,R2,R2		//R3 = -2147483648 
mem[5-1]=32'b1110_00_0_0101_0_0000_0100_000000000000; //ADC		R4 ,R0,R0		//R4 = 41
mem[6-1]=32'b1110_00_0_0010_0_0100_0101_000100000100; //SUB		R5 ,R4,R4,LSL #2	//R5 = -123
mem[7-1]=32'b1110_00_0_0110_0_0000_0110_000010100000; //SBC		R6 ,R0,R0,LSR #1	//R6 = 10
mem[8-1]=32'b1110_00_0_1100_0_0101_0111_000101000010; //ORR		R7 ,R5,R2,ASR #2	//R7 = -123
mem[9-1]=32'b1110_00_0_0000_0_0111_1000_000000000011; //AND		R8 ,R7,R3		//R8 = -2147483648
mem[10-1]=32'b1110_00_0_1111_0_0000_1001_000000000110; //MVN		R9 ,R6		//R9 = -11
mem[11-1]=32'b1110_00_0_0001_0_0100_1010_000000000101; //EOR		R10,R4,R5	//R10 = -84
mem[12-1]=32'b1110_00_0_1010_1_1000_0000_000000000110; //CMP		R8 ,R6		
mem[13-1]=32'b0001_00_0_0100_0_0001_0001_000000000001; //ADDNE		R1 ,R1,R1		//R1 = 8192
mem[14-1]=32'b1110_00_0_1000_1_1001_0000_000000001000; //TST		R9 ,R8		
mem[15-1]=32'b0000_00_0_0100_0_0010_0010_000000000010; //ADDEQ		R2 ,R2,R2   	//R2 = -1073741824
mem[16-1]=32'b1110_00_1_1101_0_0000_0000_101100000001; //MOV		R0 ,#1024		//R0 = 1024
mem[17-1]=32'b1110_01_0_0100_0_0000_0001_000000000000; //STR		R1 ,[R0],#0	//MEM[1024] = 8192
mem[18-1]=32'b1110_01_0_0100_1_0000_1011_000000000000; //LDR		R11,[R0],#0	//R11 = 8192
mem[19-1]=32'b1110_01_0_0100_0_0000_0010_000000000100; //STR		R2 ,[R0],#4	//MEM[1028] = -1073741824
mem[20-1]=32'b1110_01_0_0100_0_0000_0011_000000001000; //STR		R3 ,[R0],#8	//MEM[1032] = -2147483648
mem[21-1]=32'b1110_01_0_0100_0_0000_0100_000000001101; //STR		R4 ,[R0],#13	//MEM[1036] = 41
mem[22-1]=32'b1110_01_0_0100_0_0000_0101_000000010000; //STR		R5 ,[R0],#16	//MEM[1040] = -123
mem[23-1]=32'b1110_01_0_0100_0_0000_0110_000000010100; //STR		R6 ,[R0],#20	//MEM[1044] = 10
mem[24-1]=32'b1110_01_0_0100_1_0000_1010_000000000100; //LDR		R10,[R0],#4	//R10 = -1073741824
mem[25-1]=32'b1110_01_0_0100_0_0000_0111_000000011000; //STR		R7 ,[R0],#24	//MEM[1048] = -123
mem[26-1]=32'b1110_00_1_1101_0_0000_0001_000000000100; //MOV		R1 ,#4		//R1 = 4
mem[27-1]=32'b1110_00_1_1101_0_0000_0010_000000000000; //MOV		R2 ,#0		//R2 = 0
mem[28-1]=32'b1110_00_1_1101_0_0000_0011_000000000000; //MOV		R3 ,#0		//R3 = 0
mem[29-1]=32'b1110_00_0_0100_0_0000_0100_000100000011; //ADD		R4 ,R0,R3,LSL #2	
mem[30-1]=32'b1110_01_0_0100_1_0100_0101_000000000000; //LDR		R5 ,[R4],#0
mem[31-1]=32'b1110_01_0_0100_1_0100_0110_000000000100; //LDR		R6 ,[R4],#4
mem[32-1]=32'b1110_00_0_1010_1_0101_0000_000000000110; //CMP		R5 ,R6
mem[33-1]=32'b1100_01_0_0100_0_0100_0110_000000000000; //STRGT		R6 ,[R4],#0
mem[34-1]=32'b1100_01_0_0100_0_0100_0101_000000000100; //STRGT		R5 ,[R4],#4
mem[35-1]=32'b1110_00_1_0100_0_0011_0011_000000000001; //ADD		R3 ,R3,#1
mem[36-1]=32'b1110_00_1_1010_1_0011_0000_000000000011; //CMP		R3 ,#3
mem[37-1]=32'b1011_10_1_0_111111111111111111110111      ; //BLT		#-9
mem[38-1]=32'b1110_00_1_0100_0_0010_0010_000000000001; //ADD		R2 ,R2,#1
mem[39-1]=32'b1110_00_0_1010_1_0010_0000_000000000001; //CMP		R2 ,R1
mem[40-1]=32'b1011_10_1_0_111111111111111111110011      ; //BLT		#-13
mem[41-1]=32'b1110_01_0_0100_1_0000_0001_000000000000; //LDR		R1 ,[R0],#0	//R1 = -2147483648
mem[42-1]=32'b1110_01_0_0100_1_0000_0010_000000000100; //LDR		R2 ,[R0],#4	//R2 = -1073741824
mem[43-1]=32'b1110_01_0_0100_1_0000_0011_000000001000; //LDR		R3 ,[R0],#8	//R3 = 41
mem[44-1]=32'b1110_01_0_0100_1_0000_0100_000000001100; //LDR		R4 ,[R0],#12	//R4 = 8192
mem[45-1]=32'b1110_01_0_0100_1_0000_0101_000000010000; //LDR		R5 ,[R0],#16	//R5 = -123
mem[46-1]=32'b1110_01_0_0100_1_0000_0110_000000010100; //LDR		R6 ,[R0],#20	//R4 = 10
mem[47-1]=32'b1110_10_1_0_111111111111111111111111      ; //B		#-1
mem[48-1]=32'd0;
mem[49-1]=32'd0;
mem[50-1]=32'd0;
mem[51-1]=32'd0;
end

always @(Address) begin
    inst<=mem[Address[31:2]];
end
endmodule